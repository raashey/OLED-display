library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity character_ROM is
port (CLK : in std_logic;
      EN : in std_logic;
      ADDR : in std_logic_vector(6 downto 0);
      DATA : out std_logic_vector(7 downto 0) := "00000000");
end character_ROM;

architecture syn of character_ROM is
    type rom_type is array (0 to 127) of std_logic_vector (7 downto 0);                 
    signal ROM : rom_type:= (
	 
			"00000000", -- 0
			"00111110",
			"01010001",
			"01001001",
			"01000101",
			"00111110",
			"00000000",
			"00000000",
			
			"00000000", -- 1
			"00000000",
			"01000010",
			"01111111",
			"01000000",
			"00000000",
			"00000000",
			"00000000",
			
			"00000000", -- 2
			"01000010",
			"01100001",
			"01010001",
			"01001001",
			"01000110",
			"00000000",
			"00000000",
			
			"00000000", -- 3
			"00100001",
			"01000001",
			"01000101",
			"01001011",
			"00110001",
			"00000000",
			"00000000",
			
			"00000000", -- 4
			"00011000",
			"00010100",
			"00010010",
			"01111111",
			"00010000",
			"00000000",
			"00000000",
			
			"00000000", -- 5
			"00100111",
			"01000101",
			"01000101",
			"01000101",
			"00111001",
			"00000000",
			"00000000",
			
			"00000000", -- 6
			"00111100",
			"01001010",
			"01001001",
			"01001001",
			"00110000",
			"00000000",
			"00000000",
			
			"00000000", -- 7
			"00000001",
			"01110001",
			"00001001",
			"00000101",
			"00000011",
			"00000000",
			"00000000",
			
			"00000000", -- 8
			"00110110",
			"01001001",
			"01001001",
			"01001001",
			"00110110",
			"00000000",
			"00000000",
			
			"00000000", -- 9
			"00000110",
			"01001001",
			"01001001",
			"00101001",
			"00011110",
			"00000000",
			"00000000",
			
			"00000000", -- +
			"00001000",
			"00001000",
			"00111110",
			"00001000",
			"00001000",
			"00000000",
			"00000000",
			
			"00000000", -- -
			"00001000",
			"00001000",
			"00001000",
			"00001000",
			"00001000",
			"00000000",
			"00000000",
			
			"00000000", -- C
			"00111110",
			"01000001",
			"01000001",
			"01000001",
			"00100010",
			"00000000",
			"00000000",
			
			"00000000", -- D
			"01111111",
			"01000001",
			"01000001",
			"01000001",
			"00111110",
			"00000000",
			"00000000",
		
			"00000000", -- E
			"01111111",
			"01001001",
			"01001001",
			"01001001",
			"01000001",
			"00000000",
			"00000000",
		
			"00000000", -- F
			"01111111",
			"00001001",
			"00001001",
			"00001001",
			"00000001",
			"00000000",
			"00000000");                        

    signal rdata : std_logic_vector(7 downto 0);
begin

    rdata <= ROM(conv_integer(ADDR));

    process (CLK)
    begin
        if (CLK'event and CLK = '1') then
            if (EN = '1') then
                DATA <= rdata;
            end if;
        end if;
    end process;

end syn;
